VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO prediction
  CLASS BLOCK ;
  FOREIGN prediction ;
  ORIGIN 0.000 0.000 ;
  SIZE 965.765 BY 976.485 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 972.485 16.930 976.485 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 972.485 265.330 976.485 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 972.485 290.170 976.485 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 972.485 315.010 976.485 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 972.485 339.850 976.485 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 972.485 364.690 976.485 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 972.485 389.530 976.485 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 972.485 414.370 976.485 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 972.485 439.210 976.485 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 972.485 464.050 976.485 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 972.485 488.890 976.485 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 972.485 41.770 976.485 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 972.485 513.730 976.485 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 972.485 538.570 976.485 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 972.485 563.410 976.485 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 972.485 588.250 976.485 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 972.485 613.090 976.485 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 972.485 637.930 976.485 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 972.485 662.770 976.485 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 972.485 687.610 976.485 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 972.485 712.450 976.485 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 972.485 737.290 976.485 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 972.485 66.610 976.485 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 972.485 762.130 976.485 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 972.485 786.970 976.485 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 972.485 811.810 976.485 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 972.485 836.650 976.485 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 972.485 861.490 976.485 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 972.485 886.330 976.485 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 972.485 911.170 976.485 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 972.485 936.010 976.485 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 972.485 91.450 976.485 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 972.485 116.290 976.485 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 972.485 141.130 976.485 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 972.485 165.970 976.485 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 972.485 190.810 976.485 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 972.485 215.650 976.485 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 972.485 240.490 976.485 ;
    END
  END io_in[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 972.485 29.350 976.485 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 972.485 277.750 976.485 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 972.485 302.590 976.485 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 972.485 327.430 976.485 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 972.485 352.270 976.485 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 972.485 377.110 976.485 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 972.485 401.950 976.485 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 972.485 426.790 976.485 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 972.485 451.630 976.485 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 972.485 476.470 976.485 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 972.485 501.310 976.485 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 972.485 54.190 976.485 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 972.485 526.150 976.485 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 972.485 550.990 976.485 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 972.485 575.830 976.485 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 972.485 600.670 976.485 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 972.485 625.510 976.485 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 972.485 650.350 976.485 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 972.485 675.190 976.485 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 972.485 700.030 976.485 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 972.485 724.870 976.485 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 972.485 749.710 976.485 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 972.485 79.030 976.485 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 972.485 774.550 976.485 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 972.485 799.390 976.485 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 972.485 824.230 976.485 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 972.485 849.070 976.485 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 972.485 873.910 976.485 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 972.485 898.750 976.485 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.310 972.485 923.590 976.485 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 972.485 948.430 976.485 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 972.485 103.870 976.485 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 972.485 128.710 976.485 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 972.485 153.550 976.485 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 972.485 178.390 976.485 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 972.485 203.230 976.485 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 972.485 228.070 976.485 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 972.485 252.910 976.485 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 965.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 965.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 965.840 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wb_clk_i
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 0.000 772.710 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 0.000 801.690 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 0.000 859.650 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.330 0.000 917.610 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 0.000 946.590 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END wbs_dat_o[9]
  OBS
      LAYER nwell ;
        RECT 5.330 964.185 960.210 965.790 ;
        RECT 5.330 958.745 960.210 961.575 ;
        RECT 5.330 953.305 960.210 956.135 ;
        RECT 5.330 947.865 960.210 950.695 ;
        RECT 5.330 942.425 960.210 945.255 ;
        RECT 5.330 936.985 960.210 939.815 ;
        RECT 5.330 931.545 960.210 934.375 ;
        RECT 5.330 926.105 960.210 928.935 ;
        RECT 5.330 920.665 960.210 923.495 ;
        RECT 5.330 915.225 960.210 918.055 ;
        RECT 5.330 909.785 960.210 912.615 ;
        RECT 5.330 904.345 960.210 907.175 ;
        RECT 5.330 898.905 960.210 901.735 ;
        RECT 5.330 893.465 960.210 896.295 ;
        RECT 5.330 888.025 960.210 890.855 ;
        RECT 5.330 882.585 960.210 885.415 ;
        RECT 5.330 877.145 960.210 879.975 ;
        RECT 5.330 871.705 960.210 874.535 ;
        RECT 5.330 866.265 960.210 869.095 ;
        RECT 5.330 860.825 960.210 863.655 ;
        RECT 5.330 855.385 960.210 858.215 ;
        RECT 5.330 849.945 960.210 852.775 ;
        RECT 5.330 844.505 960.210 847.335 ;
        RECT 5.330 839.065 960.210 841.895 ;
        RECT 5.330 833.625 960.210 836.455 ;
        RECT 5.330 828.185 960.210 831.015 ;
        RECT 5.330 822.745 960.210 825.575 ;
        RECT 5.330 817.305 960.210 820.135 ;
        RECT 5.330 811.865 960.210 814.695 ;
        RECT 5.330 806.425 960.210 809.255 ;
        RECT 5.330 800.985 960.210 803.815 ;
        RECT 5.330 795.545 960.210 798.375 ;
        RECT 5.330 790.105 960.210 792.935 ;
        RECT 5.330 784.665 960.210 787.495 ;
        RECT 5.330 779.225 960.210 782.055 ;
        RECT 5.330 773.785 960.210 776.615 ;
        RECT 5.330 768.345 960.210 771.175 ;
        RECT 5.330 762.905 960.210 765.735 ;
        RECT 5.330 757.465 960.210 760.295 ;
        RECT 5.330 752.025 960.210 754.855 ;
        RECT 5.330 746.585 960.210 749.415 ;
        RECT 5.330 741.145 960.210 743.975 ;
        RECT 5.330 735.705 960.210 738.535 ;
        RECT 5.330 730.265 960.210 733.095 ;
        RECT 5.330 724.825 960.210 727.655 ;
        RECT 5.330 719.385 960.210 722.215 ;
        RECT 5.330 713.945 960.210 716.775 ;
        RECT 5.330 708.505 960.210 711.335 ;
        RECT 5.330 703.065 960.210 705.895 ;
        RECT 5.330 697.625 960.210 700.455 ;
        RECT 5.330 692.185 960.210 695.015 ;
        RECT 5.330 686.745 960.210 689.575 ;
        RECT 5.330 681.305 960.210 684.135 ;
        RECT 5.330 675.865 960.210 678.695 ;
        RECT 5.330 670.425 960.210 673.255 ;
        RECT 5.330 664.985 960.210 667.815 ;
        RECT 5.330 659.545 960.210 662.375 ;
        RECT 5.330 654.105 960.210 656.935 ;
        RECT 5.330 648.665 960.210 651.495 ;
        RECT 5.330 643.225 960.210 646.055 ;
        RECT 5.330 637.785 960.210 640.615 ;
        RECT 5.330 632.345 960.210 635.175 ;
        RECT 5.330 626.905 960.210 629.735 ;
        RECT 5.330 621.465 960.210 624.295 ;
        RECT 5.330 616.025 960.210 618.855 ;
        RECT 5.330 610.585 960.210 613.415 ;
        RECT 5.330 605.145 960.210 607.975 ;
        RECT 5.330 599.705 960.210 602.535 ;
        RECT 5.330 594.265 960.210 597.095 ;
        RECT 5.330 588.825 960.210 591.655 ;
        RECT 5.330 583.385 960.210 586.215 ;
        RECT 5.330 577.945 960.210 580.775 ;
        RECT 5.330 572.505 960.210 575.335 ;
        RECT 5.330 567.065 960.210 569.895 ;
        RECT 5.330 561.625 960.210 564.455 ;
        RECT 5.330 556.185 960.210 559.015 ;
        RECT 5.330 550.745 960.210 553.575 ;
        RECT 5.330 545.305 960.210 548.135 ;
        RECT 5.330 539.865 960.210 542.695 ;
        RECT 5.330 534.425 960.210 537.255 ;
        RECT 5.330 528.985 960.210 531.815 ;
        RECT 5.330 523.545 960.210 526.375 ;
        RECT 5.330 518.105 960.210 520.935 ;
        RECT 5.330 512.665 960.210 515.495 ;
        RECT 5.330 507.225 960.210 510.055 ;
        RECT 5.330 501.785 960.210 504.615 ;
        RECT 5.330 496.345 960.210 499.175 ;
        RECT 5.330 490.905 960.210 493.735 ;
        RECT 5.330 485.465 960.210 488.295 ;
        RECT 5.330 480.025 960.210 482.855 ;
        RECT 5.330 474.585 960.210 477.415 ;
        RECT 5.330 469.145 960.210 471.975 ;
        RECT 5.330 463.705 960.210 466.535 ;
        RECT 5.330 458.265 960.210 461.095 ;
        RECT 5.330 452.825 960.210 455.655 ;
        RECT 5.330 447.385 960.210 450.215 ;
        RECT 5.330 441.945 960.210 444.775 ;
        RECT 5.330 436.505 960.210 439.335 ;
        RECT 5.330 431.065 960.210 433.895 ;
        RECT 5.330 425.625 960.210 428.455 ;
        RECT 5.330 420.185 960.210 423.015 ;
        RECT 5.330 414.745 960.210 417.575 ;
        RECT 5.330 409.305 960.210 412.135 ;
        RECT 5.330 403.865 960.210 406.695 ;
        RECT 5.330 398.425 960.210 401.255 ;
        RECT 5.330 392.985 960.210 395.815 ;
        RECT 5.330 387.545 960.210 390.375 ;
        RECT 5.330 382.105 960.210 384.935 ;
        RECT 5.330 376.665 960.210 379.495 ;
        RECT 5.330 371.225 960.210 374.055 ;
        RECT 5.330 365.785 960.210 368.615 ;
        RECT 5.330 360.345 960.210 363.175 ;
        RECT 5.330 354.905 960.210 357.735 ;
        RECT 5.330 349.465 960.210 352.295 ;
        RECT 5.330 344.025 960.210 346.855 ;
        RECT 5.330 338.585 960.210 341.415 ;
        RECT 5.330 333.145 960.210 335.975 ;
        RECT 5.330 327.705 960.210 330.535 ;
        RECT 5.330 322.265 960.210 325.095 ;
        RECT 5.330 316.825 960.210 319.655 ;
        RECT 5.330 311.385 960.210 314.215 ;
        RECT 5.330 305.945 960.210 308.775 ;
        RECT 5.330 300.505 960.210 303.335 ;
        RECT 5.330 295.065 960.210 297.895 ;
        RECT 5.330 289.625 960.210 292.455 ;
        RECT 5.330 284.185 960.210 287.015 ;
        RECT 5.330 278.745 960.210 281.575 ;
        RECT 5.330 273.305 960.210 276.135 ;
        RECT 5.330 267.865 960.210 270.695 ;
        RECT 5.330 262.425 960.210 265.255 ;
        RECT 5.330 256.985 960.210 259.815 ;
        RECT 5.330 251.545 960.210 254.375 ;
        RECT 5.330 246.105 960.210 248.935 ;
        RECT 5.330 240.665 960.210 243.495 ;
        RECT 5.330 235.225 960.210 238.055 ;
        RECT 5.330 229.785 960.210 232.615 ;
        RECT 5.330 224.345 960.210 227.175 ;
        RECT 5.330 218.905 960.210 221.735 ;
        RECT 5.330 213.465 960.210 216.295 ;
        RECT 5.330 208.025 960.210 210.855 ;
        RECT 5.330 202.585 960.210 205.415 ;
        RECT 5.330 197.145 960.210 199.975 ;
        RECT 5.330 191.705 960.210 194.535 ;
        RECT 5.330 186.265 960.210 189.095 ;
        RECT 5.330 180.825 960.210 183.655 ;
        RECT 5.330 175.385 960.210 178.215 ;
        RECT 5.330 169.945 960.210 172.775 ;
        RECT 5.330 164.505 960.210 167.335 ;
        RECT 5.330 159.065 960.210 161.895 ;
        RECT 5.330 153.625 960.210 156.455 ;
        RECT 5.330 148.185 960.210 151.015 ;
        RECT 5.330 142.745 960.210 145.575 ;
        RECT 5.330 137.305 960.210 140.135 ;
        RECT 5.330 131.865 960.210 134.695 ;
        RECT 5.330 126.425 960.210 129.255 ;
        RECT 5.330 120.985 960.210 123.815 ;
        RECT 5.330 115.545 960.210 118.375 ;
        RECT 5.330 110.105 960.210 112.935 ;
        RECT 5.330 104.665 960.210 107.495 ;
        RECT 5.330 99.225 960.210 102.055 ;
        RECT 5.330 93.785 960.210 96.615 ;
        RECT 5.330 88.345 960.210 91.175 ;
        RECT 5.330 82.905 960.210 85.735 ;
        RECT 5.330 77.465 960.210 80.295 ;
        RECT 5.330 72.025 960.210 74.855 ;
        RECT 5.330 66.585 960.210 69.415 ;
        RECT 5.330 61.145 960.210 63.975 ;
        RECT 5.330 55.705 960.210 58.535 ;
        RECT 5.330 50.265 960.210 53.095 ;
        RECT 5.330 44.825 960.210 47.655 ;
        RECT 5.330 39.385 960.210 42.215 ;
        RECT 5.330 33.945 960.210 36.775 ;
        RECT 5.330 28.505 960.210 31.335 ;
        RECT 5.330 23.065 960.210 25.895 ;
        RECT 5.330 17.625 960.210 20.455 ;
        RECT 5.330 12.185 960.210 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 960.020 965.685 ;
      LAYER met1 ;
        RECT 5.520 10.640 961.330 970.320 ;
      LAYER met2 ;
        RECT 13.890 972.205 16.370 972.810 ;
        RECT 17.210 972.205 28.790 972.810 ;
        RECT 29.630 972.205 41.210 972.810 ;
        RECT 42.050 972.205 53.630 972.810 ;
        RECT 54.470 972.205 66.050 972.810 ;
        RECT 66.890 972.205 78.470 972.810 ;
        RECT 79.310 972.205 90.890 972.810 ;
        RECT 91.730 972.205 103.310 972.810 ;
        RECT 104.150 972.205 115.730 972.810 ;
        RECT 116.570 972.205 128.150 972.810 ;
        RECT 128.990 972.205 140.570 972.810 ;
        RECT 141.410 972.205 152.990 972.810 ;
        RECT 153.830 972.205 165.410 972.810 ;
        RECT 166.250 972.205 177.830 972.810 ;
        RECT 178.670 972.205 190.250 972.810 ;
        RECT 191.090 972.205 202.670 972.810 ;
        RECT 203.510 972.205 215.090 972.810 ;
        RECT 215.930 972.205 227.510 972.810 ;
        RECT 228.350 972.205 239.930 972.810 ;
        RECT 240.770 972.205 252.350 972.810 ;
        RECT 253.190 972.205 264.770 972.810 ;
        RECT 265.610 972.205 277.190 972.810 ;
        RECT 278.030 972.205 289.610 972.810 ;
        RECT 290.450 972.205 302.030 972.810 ;
        RECT 302.870 972.205 314.450 972.810 ;
        RECT 315.290 972.205 326.870 972.810 ;
        RECT 327.710 972.205 339.290 972.810 ;
        RECT 340.130 972.205 351.710 972.810 ;
        RECT 352.550 972.205 364.130 972.810 ;
        RECT 364.970 972.205 376.550 972.810 ;
        RECT 377.390 972.205 388.970 972.810 ;
        RECT 389.810 972.205 401.390 972.810 ;
        RECT 402.230 972.205 413.810 972.810 ;
        RECT 414.650 972.205 426.230 972.810 ;
        RECT 427.070 972.205 438.650 972.810 ;
        RECT 439.490 972.205 451.070 972.810 ;
        RECT 451.910 972.205 463.490 972.810 ;
        RECT 464.330 972.205 475.910 972.810 ;
        RECT 476.750 972.205 488.330 972.810 ;
        RECT 489.170 972.205 500.750 972.810 ;
        RECT 501.590 972.205 513.170 972.810 ;
        RECT 514.010 972.205 525.590 972.810 ;
        RECT 526.430 972.205 538.010 972.810 ;
        RECT 538.850 972.205 550.430 972.810 ;
        RECT 551.270 972.205 562.850 972.810 ;
        RECT 563.690 972.205 575.270 972.810 ;
        RECT 576.110 972.205 587.690 972.810 ;
        RECT 588.530 972.205 600.110 972.810 ;
        RECT 600.950 972.205 612.530 972.810 ;
        RECT 613.370 972.205 624.950 972.810 ;
        RECT 625.790 972.205 637.370 972.810 ;
        RECT 638.210 972.205 649.790 972.810 ;
        RECT 650.630 972.205 662.210 972.810 ;
        RECT 663.050 972.205 674.630 972.810 ;
        RECT 675.470 972.205 687.050 972.810 ;
        RECT 687.890 972.205 699.470 972.810 ;
        RECT 700.310 972.205 711.890 972.810 ;
        RECT 712.730 972.205 724.310 972.810 ;
        RECT 725.150 972.205 736.730 972.810 ;
        RECT 737.570 972.205 749.150 972.810 ;
        RECT 749.990 972.205 761.570 972.810 ;
        RECT 762.410 972.205 773.990 972.810 ;
        RECT 774.830 972.205 786.410 972.810 ;
        RECT 787.250 972.205 798.830 972.810 ;
        RECT 799.670 972.205 811.250 972.810 ;
        RECT 812.090 972.205 823.670 972.810 ;
        RECT 824.510 972.205 836.090 972.810 ;
        RECT 836.930 972.205 848.510 972.810 ;
        RECT 849.350 972.205 860.930 972.810 ;
        RECT 861.770 972.205 873.350 972.810 ;
        RECT 874.190 972.205 885.770 972.810 ;
        RECT 886.610 972.205 898.190 972.810 ;
        RECT 899.030 972.205 910.610 972.810 ;
        RECT 911.450 972.205 923.030 972.810 ;
        RECT 923.870 972.205 935.450 972.810 ;
        RECT 936.290 972.205 947.870 972.810 ;
        RECT 948.710 972.205 961.310 972.810 ;
        RECT 13.890 4.280 961.310 972.205 ;
        RECT 13.890 3.670 18.670 4.280 ;
        RECT 19.510 3.670 47.650 4.280 ;
        RECT 48.490 3.670 76.630 4.280 ;
        RECT 77.470 3.670 105.610 4.280 ;
        RECT 106.450 3.670 134.590 4.280 ;
        RECT 135.430 3.670 163.570 4.280 ;
        RECT 164.410 3.670 192.550 4.280 ;
        RECT 193.390 3.670 221.530 4.280 ;
        RECT 222.370 3.670 250.510 4.280 ;
        RECT 251.350 3.670 279.490 4.280 ;
        RECT 280.330 3.670 308.470 4.280 ;
        RECT 309.310 3.670 337.450 4.280 ;
        RECT 338.290 3.670 366.430 4.280 ;
        RECT 367.270 3.670 395.410 4.280 ;
        RECT 396.250 3.670 424.390 4.280 ;
        RECT 425.230 3.670 453.370 4.280 ;
        RECT 454.210 3.670 482.350 4.280 ;
        RECT 483.190 3.670 511.330 4.280 ;
        RECT 512.170 3.670 540.310 4.280 ;
        RECT 541.150 3.670 569.290 4.280 ;
        RECT 570.130 3.670 598.270 4.280 ;
        RECT 599.110 3.670 627.250 4.280 ;
        RECT 628.090 3.670 656.230 4.280 ;
        RECT 657.070 3.670 685.210 4.280 ;
        RECT 686.050 3.670 714.190 4.280 ;
        RECT 715.030 3.670 743.170 4.280 ;
        RECT 744.010 3.670 772.150 4.280 ;
        RECT 772.990 3.670 801.130 4.280 ;
        RECT 801.970 3.670 830.110 4.280 ;
        RECT 830.950 3.670 859.090 4.280 ;
        RECT 859.930 3.670 888.070 4.280 ;
        RECT 888.910 3.670 917.050 4.280 ;
        RECT 917.890 3.670 946.030 4.280 ;
        RECT 946.870 3.670 961.310 4.280 ;
      LAYER met3 ;
        RECT 13.865 10.715 961.335 972.220 ;
      LAYER met4 ;
        RECT 85.855 966.240 948.225 972.225 ;
        RECT 85.855 115.775 97.440 966.240 ;
        RECT 99.840 115.775 174.240 966.240 ;
        RECT 176.640 115.775 251.040 966.240 ;
        RECT 253.440 115.775 327.840 966.240 ;
        RECT 330.240 115.775 404.640 966.240 ;
        RECT 407.040 115.775 481.440 966.240 ;
        RECT 483.840 115.775 558.240 966.240 ;
        RECT 560.640 115.775 635.040 966.240 ;
        RECT 637.440 115.775 711.840 966.240 ;
        RECT 714.240 115.775 788.640 966.240 ;
        RECT 791.040 115.775 865.440 966.240 ;
        RECT 867.840 115.775 942.240 966.240 ;
        RECT 944.640 115.775 948.225 966.240 ;
  END
END prediction
END LIBRARY

