magic
tech sky130B
magscale 1 2
timestamp 1658125919
<< nwell >>
rect 1066 192837 192042 193158
rect 1066 191749 192042 192315
rect 1066 190661 192042 191227
rect 1066 189573 192042 190139
rect 1066 188485 192042 189051
rect 1066 187397 192042 187963
rect 1066 186309 192042 186875
rect 1066 185221 192042 185787
rect 1066 184133 192042 184699
rect 1066 183045 192042 183611
rect 1066 181957 192042 182523
rect 1066 180869 192042 181435
rect 1066 179781 192042 180347
rect 1066 178693 192042 179259
rect 1066 177605 192042 178171
rect 1066 176517 192042 177083
rect 1066 175429 192042 175995
rect 1066 174341 192042 174907
rect 1066 173253 192042 173819
rect 1066 172165 192042 172731
rect 1066 171077 192042 171643
rect 1066 169989 192042 170555
rect 1066 168901 192042 169467
rect 1066 167813 192042 168379
rect 1066 166725 192042 167291
rect 1066 165637 192042 166203
rect 1066 164549 192042 165115
rect 1066 163461 192042 164027
rect 1066 162373 192042 162939
rect 1066 161285 192042 161851
rect 1066 160197 192042 160763
rect 1066 159109 192042 159675
rect 1066 158021 192042 158587
rect 1066 156933 192042 157499
rect 1066 155845 192042 156411
rect 1066 154757 192042 155323
rect 1066 153669 192042 154235
rect 1066 152581 192042 153147
rect 1066 151493 192042 152059
rect 1066 150405 192042 150971
rect 1066 149317 192042 149883
rect 1066 148229 192042 148795
rect 1066 147141 192042 147707
rect 1066 146053 192042 146619
rect 1066 144965 192042 145531
rect 1066 143877 192042 144443
rect 1066 142789 192042 143355
rect 1066 141701 192042 142267
rect 1066 140613 192042 141179
rect 1066 139525 192042 140091
rect 1066 138437 192042 139003
rect 1066 137349 192042 137915
rect 1066 136261 192042 136827
rect 1066 135173 192042 135739
rect 1066 134085 192042 134651
rect 1066 132997 192042 133563
rect 1066 131909 192042 132475
rect 1066 130821 192042 131387
rect 1066 129733 192042 130299
rect 1066 128645 192042 129211
rect 1066 127557 192042 128123
rect 1066 126469 192042 127035
rect 1066 125381 192042 125947
rect 1066 124293 192042 124859
rect 1066 123205 192042 123771
rect 1066 122117 192042 122683
rect 1066 121029 192042 121595
rect 1066 119941 192042 120507
rect 1066 118853 192042 119419
rect 1066 117765 192042 118331
rect 1066 116677 192042 117243
rect 1066 115589 192042 116155
rect 1066 114501 192042 115067
rect 1066 113413 192042 113979
rect 1066 112325 192042 112891
rect 1066 111237 192042 111803
rect 1066 110149 192042 110715
rect 1066 109061 192042 109627
rect 1066 107973 192042 108539
rect 1066 106885 192042 107451
rect 1066 105797 192042 106363
rect 1066 104709 192042 105275
rect 1066 103621 192042 104187
rect 1066 102533 192042 103099
rect 1066 101445 192042 102011
rect 1066 100357 192042 100923
rect 1066 99269 192042 99835
rect 1066 98181 192042 98747
rect 1066 97093 192042 97659
rect 1066 96005 192042 96571
rect 1066 94917 192042 95483
rect 1066 93829 192042 94395
rect 1066 92741 192042 93307
rect 1066 91653 192042 92219
rect 1066 90565 192042 91131
rect 1066 89477 192042 90043
rect 1066 88389 192042 88955
rect 1066 87301 192042 87867
rect 1066 86213 192042 86779
rect 1066 85125 192042 85691
rect 1066 84037 192042 84603
rect 1066 82949 192042 83515
rect 1066 81861 192042 82427
rect 1066 80773 192042 81339
rect 1066 79685 192042 80251
rect 1066 78597 192042 79163
rect 1066 77509 192042 78075
rect 1066 76421 192042 76987
rect 1066 75333 192042 75899
rect 1066 74245 192042 74811
rect 1066 73157 192042 73723
rect 1066 72069 192042 72635
rect 1066 70981 192042 71547
rect 1066 69893 192042 70459
rect 1066 68805 192042 69371
rect 1066 67717 192042 68283
rect 1066 66629 192042 67195
rect 1066 65541 192042 66107
rect 1066 64453 192042 65019
rect 1066 63365 192042 63931
rect 1066 62277 192042 62843
rect 1066 61189 192042 61755
rect 1066 60101 192042 60667
rect 1066 59013 192042 59579
rect 1066 57925 192042 58491
rect 1066 56837 192042 57403
rect 1066 55749 192042 56315
rect 1066 54661 192042 55227
rect 1066 53573 192042 54139
rect 1066 52485 192042 53051
rect 1066 51397 192042 51963
rect 1066 50309 192042 50875
rect 1066 49221 192042 49787
rect 1066 48133 192042 48699
rect 1066 47045 192042 47611
rect 1066 45957 192042 46523
rect 1066 44869 192042 45435
rect 1066 43781 192042 44347
rect 1066 42693 192042 43259
rect 1066 41605 192042 42171
rect 1066 40517 192042 41083
rect 1066 39429 192042 39995
rect 1066 38341 192042 38907
rect 1066 37253 192042 37819
rect 1066 36165 192042 36731
rect 1066 35077 192042 35643
rect 1066 33989 192042 34555
rect 1066 32901 192042 33467
rect 1066 31813 192042 32379
rect 1066 30725 192042 31291
rect 1066 29637 192042 30203
rect 1066 28549 192042 29115
rect 1066 27461 192042 28027
rect 1066 26373 192042 26939
rect 1066 25285 192042 25851
rect 1066 24197 192042 24763
rect 1066 23109 192042 23675
rect 1066 22021 192042 22587
rect 1066 20933 192042 21499
rect 1066 19845 192042 20411
rect 1066 18757 192042 19323
rect 1066 17669 192042 18235
rect 1066 16581 192042 17147
rect 1066 15493 192042 16059
rect 1066 14405 192042 14971
rect 1066 13317 192042 13883
rect 1066 12229 192042 12795
rect 1066 11141 192042 11707
rect 1066 10053 192042 10619
rect 1066 8965 192042 9531
rect 1066 7877 192042 8443
rect 1066 6789 192042 7355
rect 1066 5701 192042 6267
rect 1066 4613 192042 5179
rect 1066 3525 192042 4091
rect 1066 2437 192042 3003
<< obsli1 >>
rect 1104 2159 192004 193137
<< obsm1 >>
rect 1104 2128 192266 194064
<< metal2 >>
rect 3330 194497 3386 195297
rect 5814 194497 5870 195297
rect 8298 194497 8354 195297
rect 10782 194497 10838 195297
rect 13266 194497 13322 195297
rect 15750 194497 15806 195297
rect 18234 194497 18290 195297
rect 20718 194497 20774 195297
rect 23202 194497 23258 195297
rect 25686 194497 25742 195297
rect 28170 194497 28226 195297
rect 30654 194497 30710 195297
rect 33138 194497 33194 195297
rect 35622 194497 35678 195297
rect 38106 194497 38162 195297
rect 40590 194497 40646 195297
rect 43074 194497 43130 195297
rect 45558 194497 45614 195297
rect 48042 194497 48098 195297
rect 50526 194497 50582 195297
rect 53010 194497 53066 195297
rect 55494 194497 55550 195297
rect 57978 194497 58034 195297
rect 60462 194497 60518 195297
rect 62946 194497 63002 195297
rect 65430 194497 65486 195297
rect 67914 194497 67970 195297
rect 70398 194497 70454 195297
rect 72882 194497 72938 195297
rect 75366 194497 75422 195297
rect 77850 194497 77906 195297
rect 80334 194497 80390 195297
rect 82818 194497 82874 195297
rect 85302 194497 85358 195297
rect 87786 194497 87842 195297
rect 90270 194497 90326 195297
rect 92754 194497 92810 195297
rect 95238 194497 95294 195297
rect 97722 194497 97778 195297
rect 100206 194497 100262 195297
rect 102690 194497 102746 195297
rect 105174 194497 105230 195297
rect 107658 194497 107714 195297
rect 110142 194497 110198 195297
rect 112626 194497 112682 195297
rect 115110 194497 115166 195297
rect 117594 194497 117650 195297
rect 120078 194497 120134 195297
rect 122562 194497 122618 195297
rect 125046 194497 125102 195297
rect 127530 194497 127586 195297
rect 130014 194497 130070 195297
rect 132498 194497 132554 195297
rect 134982 194497 135038 195297
rect 137466 194497 137522 195297
rect 139950 194497 140006 195297
rect 142434 194497 142490 195297
rect 144918 194497 144974 195297
rect 147402 194497 147458 195297
rect 149886 194497 149942 195297
rect 152370 194497 152426 195297
rect 154854 194497 154910 195297
rect 157338 194497 157394 195297
rect 159822 194497 159878 195297
rect 162306 194497 162362 195297
rect 164790 194497 164846 195297
rect 167274 194497 167330 195297
rect 169758 194497 169814 195297
rect 172242 194497 172298 195297
rect 174726 194497 174782 195297
rect 177210 194497 177266 195297
rect 179694 194497 179750 195297
rect 182178 194497 182234 195297
rect 184662 194497 184718 195297
rect 187146 194497 187202 195297
rect 189630 194497 189686 195297
rect 3790 0 3846 800
rect 9586 0 9642 800
rect 15382 0 15438 800
rect 21178 0 21234 800
rect 26974 0 27030 800
rect 32770 0 32826 800
rect 38566 0 38622 800
rect 44362 0 44418 800
rect 50158 0 50214 800
rect 55954 0 56010 800
rect 61750 0 61806 800
rect 67546 0 67602 800
rect 73342 0 73398 800
rect 79138 0 79194 800
rect 84934 0 84990 800
rect 90730 0 90786 800
rect 96526 0 96582 800
rect 102322 0 102378 800
rect 108118 0 108174 800
rect 113914 0 113970 800
rect 119710 0 119766 800
rect 125506 0 125562 800
rect 131302 0 131358 800
rect 137098 0 137154 800
rect 142894 0 142950 800
rect 148690 0 148746 800
rect 154486 0 154542 800
rect 160282 0 160338 800
rect 166078 0 166134 800
rect 171874 0 171930 800
rect 177670 0 177726 800
rect 183466 0 183522 800
rect 189262 0 189318 800
<< obsm2 >>
rect 2778 194441 3274 194562
rect 3442 194441 5758 194562
rect 5926 194441 8242 194562
rect 8410 194441 10726 194562
rect 10894 194441 13210 194562
rect 13378 194441 15694 194562
rect 15862 194441 18178 194562
rect 18346 194441 20662 194562
rect 20830 194441 23146 194562
rect 23314 194441 25630 194562
rect 25798 194441 28114 194562
rect 28282 194441 30598 194562
rect 30766 194441 33082 194562
rect 33250 194441 35566 194562
rect 35734 194441 38050 194562
rect 38218 194441 40534 194562
rect 40702 194441 43018 194562
rect 43186 194441 45502 194562
rect 45670 194441 47986 194562
rect 48154 194441 50470 194562
rect 50638 194441 52954 194562
rect 53122 194441 55438 194562
rect 55606 194441 57922 194562
rect 58090 194441 60406 194562
rect 60574 194441 62890 194562
rect 63058 194441 65374 194562
rect 65542 194441 67858 194562
rect 68026 194441 70342 194562
rect 70510 194441 72826 194562
rect 72994 194441 75310 194562
rect 75478 194441 77794 194562
rect 77962 194441 80278 194562
rect 80446 194441 82762 194562
rect 82930 194441 85246 194562
rect 85414 194441 87730 194562
rect 87898 194441 90214 194562
rect 90382 194441 92698 194562
rect 92866 194441 95182 194562
rect 95350 194441 97666 194562
rect 97834 194441 100150 194562
rect 100318 194441 102634 194562
rect 102802 194441 105118 194562
rect 105286 194441 107602 194562
rect 107770 194441 110086 194562
rect 110254 194441 112570 194562
rect 112738 194441 115054 194562
rect 115222 194441 117538 194562
rect 117706 194441 120022 194562
rect 120190 194441 122506 194562
rect 122674 194441 124990 194562
rect 125158 194441 127474 194562
rect 127642 194441 129958 194562
rect 130126 194441 132442 194562
rect 132610 194441 134926 194562
rect 135094 194441 137410 194562
rect 137578 194441 139894 194562
rect 140062 194441 142378 194562
rect 142546 194441 144862 194562
rect 145030 194441 147346 194562
rect 147514 194441 149830 194562
rect 149998 194441 152314 194562
rect 152482 194441 154798 194562
rect 154966 194441 157282 194562
rect 157450 194441 159766 194562
rect 159934 194441 162250 194562
rect 162418 194441 164734 194562
rect 164902 194441 167218 194562
rect 167386 194441 169702 194562
rect 169870 194441 172186 194562
rect 172354 194441 174670 194562
rect 174838 194441 177154 194562
rect 177322 194441 179638 194562
rect 179806 194441 182122 194562
rect 182290 194441 184606 194562
rect 184774 194441 187090 194562
rect 187258 194441 189574 194562
rect 189742 194441 192262 194562
rect 2778 856 192262 194441
rect 2778 734 3734 856
rect 3902 734 9530 856
rect 9698 734 15326 856
rect 15494 734 21122 856
rect 21290 734 26918 856
rect 27086 734 32714 856
rect 32882 734 38510 856
rect 38678 734 44306 856
rect 44474 734 50102 856
rect 50270 734 55898 856
rect 56066 734 61694 856
rect 61862 734 67490 856
rect 67658 734 73286 856
rect 73454 734 79082 856
rect 79250 734 84878 856
rect 85046 734 90674 856
rect 90842 734 96470 856
rect 96638 734 102266 856
rect 102434 734 108062 856
rect 108230 734 113858 856
rect 114026 734 119654 856
rect 119822 734 125450 856
rect 125618 734 131246 856
rect 131414 734 137042 856
rect 137210 734 142838 856
rect 143006 734 148634 856
rect 148802 734 154430 856
rect 154598 734 160226 856
rect 160394 734 166022 856
rect 166190 734 171818 856
rect 171986 734 177614 856
rect 177782 734 183410 856
rect 183578 734 189206 856
rect 189374 734 192262 856
<< obsm3 >>
rect 2773 2143 192267 194444
<< metal4 >>
rect 4208 2128 4528 193168
rect 19568 2128 19888 193168
rect 34928 2128 35248 193168
rect 50288 2128 50608 193168
rect 65648 2128 65968 193168
rect 81008 2128 81328 193168
rect 96368 2128 96688 193168
rect 111728 2128 112048 193168
rect 127088 2128 127408 193168
rect 142448 2128 142768 193168
rect 157808 2128 158128 193168
rect 173168 2128 173488 193168
rect 188528 2128 188848 193168
<< obsm4 >>
rect 17171 193248 189645 194445
rect 17171 23155 19488 193248
rect 19968 23155 34848 193248
rect 35328 23155 50208 193248
rect 50688 23155 65568 193248
rect 66048 23155 80928 193248
rect 81408 23155 96288 193248
rect 96768 23155 111648 193248
rect 112128 23155 127008 193248
rect 127488 23155 142368 193248
rect 142848 23155 157728 193248
rect 158208 23155 173088 193248
rect 173568 23155 188448 193248
rect 188928 23155 189645 193248
<< labels >>
rlabel metal2 s 3330 194497 3386 195297 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 53010 194497 53066 195297 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 57978 194497 58034 195297 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 62946 194497 63002 195297 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 67914 194497 67970 195297 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 72882 194497 72938 195297 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 77850 194497 77906 195297 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 82818 194497 82874 195297 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 87786 194497 87842 195297 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 92754 194497 92810 195297 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 97722 194497 97778 195297 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8298 194497 8354 195297 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 102690 194497 102746 195297 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 107658 194497 107714 195297 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 112626 194497 112682 195297 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 117594 194497 117650 195297 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 122562 194497 122618 195297 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 127530 194497 127586 195297 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 132498 194497 132554 195297 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 137466 194497 137522 195297 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 142434 194497 142490 195297 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 147402 194497 147458 195297 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 13266 194497 13322 195297 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 152370 194497 152426 195297 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 157338 194497 157394 195297 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 162306 194497 162362 195297 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 167274 194497 167330 195297 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 172242 194497 172298 195297 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 177210 194497 177266 195297 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 182178 194497 182234 195297 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 187146 194497 187202 195297 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 18234 194497 18290 195297 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 23202 194497 23258 195297 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 28170 194497 28226 195297 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 33138 194497 33194 195297 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 38106 194497 38162 195297 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 43074 194497 43130 195297 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 48042 194497 48098 195297 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5814 194497 5870 195297 6 io_out[0]
port 39 nsew signal output
rlabel metal2 s 55494 194497 55550 195297 6 io_out[10]
port 40 nsew signal output
rlabel metal2 s 60462 194497 60518 195297 6 io_out[11]
port 41 nsew signal output
rlabel metal2 s 65430 194497 65486 195297 6 io_out[12]
port 42 nsew signal output
rlabel metal2 s 70398 194497 70454 195297 6 io_out[13]
port 43 nsew signal output
rlabel metal2 s 75366 194497 75422 195297 6 io_out[14]
port 44 nsew signal output
rlabel metal2 s 80334 194497 80390 195297 6 io_out[15]
port 45 nsew signal output
rlabel metal2 s 85302 194497 85358 195297 6 io_out[16]
port 46 nsew signal output
rlabel metal2 s 90270 194497 90326 195297 6 io_out[17]
port 47 nsew signal output
rlabel metal2 s 95238 194497 95294 195297 6 io_out[18]
port 48 nsew signal output
rlabel metal2 s 100206 194497 100262 195297 6 io_out[19]
port 49 nsew signal output
rlabel metal2 s 10782 194497 10838 195297 6 io_out[1]
port 50 nsew signal output
rlabel metal2 s 105174 194497 105230 195297 6 io_out[20]
port 51 nsew signal output
rlabel metal2 s 110142 194497 110198 195297 6 io_out[21]
port 52 nsew signal output
rlabel metal2 s 115110 194497 115166 195297 6 io_out[22]
port 53 nsew signal output
rlabel metal2 s 120078 194497 120134 195297 6 io_out[23]
port 54 nsew signal output
rlabel metal2 s 125046 194497 125102 195297 6 io_out[24]
port 55 nsew signal output
rlabel metal2 s 130014 194497 130070 195297 6 io_out[25]
port 56 nsew signal output
rlabel metal2 s 134982 194497 135038 195297 6 io_out[26]
port 57 nsew signal output
rlabel metal2 s 139950 194497 140006 195297 6 io_out[27]
port 58 nsew signal output
rlabel metal2 s 144918 194497 144974 195297 6 io_out[28]
port 59 nsew signal output
rlabel metal2 s 149886 194497 149942 195297 6 io_out[29]
port 60 nsew signal output
rlabel metal2 s 15750 194497 15806 195297 6 io_out[2]
port 61 nsew signal output
rlabel metal2 s 154854 194497 154910 195297 6 io_out[30]
port 62 nsew signal output
rlabel metal2 s 159822 194497 159878 195297 6 io_out[31]
port 63 nsew signal output
rlabel metal2 s 164790 194497 164846 195297 6 io_out[32]
port 64 nsew signal output
rlabel metal2 s 169758 194497 169814 195297 6 io_out[33]
port 65 nsew signal output
rlabel metal2 s 174726 194497 174782 195297 6 io_out[34]
port 66 nsew signal output
rlabel metal2 s 179694 194497 179750 195297 6 io_out[35]
port 67 nsew signal output
rlabel metal2 s 184662 194497 184718 195297 6 io_out[36]
port 68 nsew signal output
rlabel metal2 s 189630 194497 189686 195297 6 io_out[37]
port 69 nsew signal output
rlabel metal2 s 20718 194497 20774 195297 6 io_out[3]
port 70 nsew signal output
rlabel metal2 s 25686 194497 25742 195297 6 io_out[4]
port 71 nsew signal output
rlabel metal2 s 30654 194497 30710 195297 6 io_out[5]
port 72 nsew signal output
rlabel metal2 s 35622 194497 35678 195297 6 io_out[6]
port 73 nsew signal output
rlabel metal2 s 40590 194497 40646 195297 6 io_out[7]
port 74 nsew signal output
rlabel metal2 s 45558 194497 45614 195297 6 io_out[8]
port 75 nsew signal output
rlabel metal2 s 50526 194497 50582 195297 6 io_out[9]
port 76 nsew signal output
rlabel metal4 s 4208 2128 4528 193168 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 193168 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 193168 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 193168 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 193168 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 193168 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 193168 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 193168 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 193168 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 193168 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 193168 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 193168 6 vssd1
port 78 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 193168 6 vssd1
port 78 nsew ground bidirectional
rlabel metal2 s 3790 0 3846 800 6 wb_clk_i
port 79 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[0]
port 80 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_o[10]
port 81 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_o[11]
port 82 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 wbs_dat_o[12]
port 83 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_o[13]
port 84 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 wbs_dat_o[14]
port 85 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 wbs_dat_o[15]
port 86 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 wbs_dat_o[16]
port 87 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 wbs_dat_o[17]
port 88 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 wbs_dat_o[18]
port 89 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 wbs_dat_o[19]
port 90 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[1]
port 91 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 wbs_dat_o[20]
port 92 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 wbs_dat_o[21]
port 93 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 wbs_dat_o[22]
port 94 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 wbs_dat_o[23]
port 95 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 wbs_dat_o[24]
port 96 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 wbs_dat_o[25]
port 97 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 wbs_dat_o[26]
port 98 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 wbs_dat_o[27]
port 99 nsew signal output
rlabel metal2 s 171874 0 171930 800 6 wbs_dat_o[28]
port 100 nsew signal output
rlabel metal2 s 177670 0 177726 800 6 wbs_dat_o[29]
port 101 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[2]
port 102 nsew signal output
rlabel metal2 s 183466 0 183522 800 6 wbs_dat_o[30]
port 103 nsew signal output
rlabel metal2 s 189262 0 189318 800 6 wbs_dat_o[31]
port 104 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[3]
port 105 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[4]
port 106 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[5]
port 107 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[6]
port 108 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_o[7]
port 109 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_o[8]
port 110 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_o[9]
port 111 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 193153 195297
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 99348178
string GDS_FILE /home/bn/mpw7_test/openlane/prediction/runs/22_07_18_16_45/results/signoff/prediction.magic.gds
string GDS_START 1656610
<< end >>

